---------------------------------------------------------------------------
--
--  Title: Hardware Thread User Logic Quicksort
--  Thread implements the quicksort algorithm
--  Passed in argument is a pointer to following struct
-- struct sortData {
--   int * startData; //pointer to start of array
--   int * endData; //pointer to end of array
--   int cacheOption // 1 operate on data where it is, 0 copy into HWTI first
--  There is not return argument, the HWT just sorts the data.
--
---------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_misc.all;

library Unisim;
use Unisim.all;

---------------------------------------------------------------------------
-- Port declarations
---------------------------------------------------------------------------
-- Definition of Ports:
--
--  Misc. Signals
--    clock
--
--  HWTI to HWTUL interconnect
--    intrfc2thrd_address      32 bits   memory    
--    intrfc2thrd_value        32 bits   memory    function
--    intrfc2thrd_function     16 bits                       control
--    intrfc2thrd_goWait        1 bits                       control
--
--  HWTUL to HWTI interconnect
--    thrd2intrfc_address      32 bits   memory
--    thrd2intrfc_value        32 bits   memory    function
--    thrd2intrfc_function     16 bits             function
--    thrd2intrfc_opcode        6 bits   memory    function
--

---------------------------------------------------------------------------
-- Thread Manager Entity section
---------------------------------------------------------------------------

entity user_logic_hwtul is
  port (
    clock : in std_logic;
    intrfc2thrd_address : in std_logic_vector(0 to 31);
    intrfc2thrd_value : in std_logic_vector(0 to 31);
    intrfc2thrd_function : in std_logic_vector(0 to 15);
    intrfc2thrd_goWait : in std_logic;

    thrd2intrfc_address : out std_logic_vector(0 to 31);
    thrd2intrfc_value : out std_logic_vector(0 to 31);
    thrd2intrfc_function : out std_logic_vector(0 to 15);
    thrd2intrfc_opcode : out std_logic_vector(0 to 5)
  );
end entity user_logic_hwtul;

---------------------------------------------------------------------------
-- Architecture section
---------------------------------------------------------------------------

architecture IMP of user_logic_hwtul is

---------------------------------------------------------------------------
-- Signal declarations
---------------------------------------------------------------------------

  type state_machine is (
    FUNCTION_RESET,
    FUNCTION_USER_SELECT,
    FUNCTION_START,
	READ_ARGS_1,
	READ_ARGS_2,
	READ_ARGS_3,
	READ_ARGS_4,
	READ_ARGS_5,
	FORLOOP_1,
	FORLOOP_2,
	FORLOOP_3,
	FORLOOP_4,
	WHILE_A_1,
	WHILE_A_2,
	WHILE_A_3,
	WHILE_B_1,
	WHILE_B_2,
	WHILE_B_3,
	WHILE_B_4,
	WHILE_B_5,
	WHILE_B_6,
	FLUSH_1,
	FLUSH_2,
    EXIT_THREAD,
    EXIT_THREAD_1,
    WAIT_STATE,
    ERROR_STATE);

  -- Function definitions
  constant U_FUNCTION_RESET                    : std_logic_vector(0 to 15) := x"0000";
  constant U_FUNCTION_WAIT                     : std_logic_vector(0 to 15) := x"0001";
  constant U_FUNCTION_USER_SELECT              : std_logic_vector(0 to 15) := x"0002";
  constant U_FUNCTION_START                    : std_logic_vector(0 to 15) := x"0003";

  -- Range 0003 to 7999 reserved for user logic's state machine
  -- Range 8000 to 9999 reserved for system calls
  constant FUNCTION_HTHREAD_ATTR_INIT          : std_logic_vector(0 to 15) := x"8000";
  constant FUNCTION_HTHREAD_ATTR_DESTROY       : std_logic_vector(0 to 15) := x"8001";
  constant FUNCTION_HTHREAD_CREATE             : std_logic_vector(0 to 15) := x"8010";
  constant FUNCTION_HTHREAD_JOIN               : std_logic_vector(0 to 15) := x"8011";
  constant FUNCTION_HTHREAD_SELF               : std_logic_vector(0 to 15) := x"8012";
  constant FUNCTION_HTHREAD_YIELD              : std_logic_vector(0 to 15) := x"8013";
  constant FUNCTION_HTHREAD_EQUAL              : std_logic_vector(0 to 15) := x"8014";
  constant FUNCTION_HTHREAD_EXIT               : std_logic_vector(0 to 15) := x"8015";
  constant FUNCTION_HTHREAD_EXIT_ERROR         : std_logic_vector(0 to 15) := x"8016";
  constant FUNCTION_HTHREAD_MUTEXATTR_INIT     : std_logic_vector(0 to 15) := x"8020";
  constant FUNCTION_HTHREAD_MUTEXATTR_DESTROY  : std_logic_vector(0 to 15) := x"8021";
  constant FUNCTION_HTHREAD_MUTEXATTR_SETNUM   : std_logic_vector(0 to 15) := x"8022";
  constant FUNCTION_HTHREAD_MUTEXATTR_GETNUM   : std_logic_vector(0 to 15) := x"8023";
  constant FUNCTION_HTHREAD_MUTEX_INIT         : std_logic_vector(0 to 15) := x"8030";
  constant FUNCTION_HTHREAD_MUTEX_DESTROY      : std_logic_vector(0 to 15) := x"8031";
  constant FUNCTION_HTHREAD_MUTEX_LOCK         : std_logic_vector(0 to 15) := x"8032";
  constant FUNCTION_HTHREAD_MUTEX_UNLOCK       : std_logic_vector(0 to 15) := x"8033";
  constant FUNCTION_HTHREAD_MUTEX_TRYLOCK      : std_logic_vector(0 to 15) := x"8034";
  constant FUNCTION_HTHREAD_CONDATTR_INIT      : std_logic_vector(0 to 15) := x"8040";
  constant FUNCTION_HTHREAD_CONDATTR_DESTROY   : std_logic_vector(0 to 15) := x"8041";
  constant FUNCTION_HTHREAD_CONDATTR_SETNUM    : std_logic_vector(0 to 15) := x"8042";
  constant FUNCTION_HTHREAD_CONDATTR_GETNUM    : std_logic_vector(0 to 15) := x"8043";
  constant FUNCTION_HTHREAD_COND_INIT          : std_logic_vector(0 to 15) := x"8050";
  constant FUNCTION_HTHREAD_COND_DESTROY       : std_logic_vector(0 to 15) := x"8051";
  constant FUNCTION_HTHREAD_COND_SIGNAL        : std_logic_vector(0 to 15) := x"8052";
  constant FUNCTION_HTHREAD_COND_BROADCAST     : std_logic_vector(0 to 15) := x"8053";
  constant FUNCTION_HTHREAD_COND_WAIT          : std_logic_vector(0 to 15) := x"8054";
  -- Ranged A000 to FFFF reserved for supported library calls
  constant FUNCTION_MALLOC                     : std_logic_vector(0 to 15) := x"A000";
  constant FUNCTION_CALLOC                     : std_logic_vector(0 to 15) := x"A001";
  constant FUNCTION_FREE                       : std_logic_vector(0 to 15) := x"A002";
  constant FUNCTION_MEMCPY                     : std_logic_vector(0 to 15) := x"A100";

  -- user_opcode Constants
  constant OPCODE_NOOP                         : std_logic_vector(0 to 5) := "000000";
  -- Memory sub-interface specific opcodes
  constant OPCODE_LOAD                         : std_logic_vector(0 to 5) := "000001";
  constant OPCODE_STORE                        : std_logic_vector(0 to 5) := "000010";
  constant OPCODE_DECLARE                      : std_logic_vector(0 to 5) := "000011";
  constant OPCODE_READ                         : std_logic_vector(0 to 5) := "000100";
  constant OPCODE_WRITE                        : std_logic_vector(0 to 5) := "000101";
  constant OPCODE_ADDRESS                      : std_logic_vector(0 to 5) := "000110";
  -- Function sub-interface specific opcodes
  constant OPCODE_PUSH                         : std_logic_vector(0 to 5) := "010000";
  constant OPCODE_POP                          : std_logic_vector(0 to 5) := "010001";
  constant OPCODE_CALL                         : std_logic_vector(0 to 5) := "010010";
  constant OPCODE_RETURN                       : std_logic_vector(0 to 5) := "010011";

  constant Z32 : std_logic_vector(0 to 31) := (others => '0');

  constant MAX_SIZE : std_logic_vector(0 to 31) := x"00000400";

  signal current_state, next_state : state_machine := FUNCTION_RESET;
  signal return_state, return_state_next : state_machine := FUNCTION_RESET;
  signal arg, arg_next : std_logic_vector(0 to 31);
  signal bufer, buffer_next : std_logic_vector(0 to 31);
  signal bufLen, bufLen_next : std_logic_vector(0 to 31);
  signal outputIndex, outputIndex_next : std_logic_vector(0 to 31);
  signal index, index_next : std_logic_vector(0 to 31);
  signal len, len_next : std_logic_vector(0 to 31);
  signal pos, pos_next : std_logic_vector(0 to 31);
  signal inputData, inputData_next : std_logic_vector(0 to 31);
  signal outputData, outputData_next : std_logic_vector(0 to 31);
  signal count, count_next : std_logic_vector(0 to 31);

  signal toUser_address : std_logic_vector(0 to 31);
  signal toUser_value : std_logic_vector(0 to 31);
  signal toUser_function : std_logic_vector(0 to 15);
  signal toUser_goWait : std_logic;

---------------------------------------------------------------------------
-- Begin architecture
---------------------------------------------------------------------------

begin -- architecture IMP

  HWTUL_STATE_PROCESS : process (clock) is
  begin
    
    if (clock'event and (clock = '1')) then
      toUser_address <= intrfc2thrd_address;
      toUser_value <= intrfc2thrd_value;
      toUser_function <= intrfc2thrd_function;
      toUser_goWait <= intrfc2thrd_goWait;

	  arg <= arg_next;
	  bufer <= buffer_next;
	  bufLen <= bufLen_next;
	  outputIndex <= outputIndex_next;
	  index <= index_next;
	  len <= len_next;
	  pos <= pos_next;
	  inputData <= inputData_next;
	  outputData <= outputData_next;
	  count <= count_next;
      return_state <= return_state_next;

      -- Find out if the HWTI is tell us what to do
      if (intrfc2thrd_goWait = '1') then
        case intrfc2thrd_function is
          -- Typically the HWTI will tell us to control our own destiny
          when U_FUNCTION_USER_SELECT =>
            current_state <= next_state;

          -- List all the functions the HWTI could tell us to run
          when U_FUNCTION_RESET =>
            current_state <= FUNCTION_RESET;
          when U_FUNCTION_START =>
            current_state <= FUNCTION_START;

          -- If the HWTI tells us to do something we don't know, error
          when OTHERS =>
            current_state <= ERROR_STATE;
        end case;
      else
        current_state <= WAIT_STATE;
      end if;
    end if;
  end process HWTUL_STATE_PROCESS;


  HWTUL_STATE_MACHINE : process (current_state) is
  begin

    -- Default register assignments
    thrd2intrfc_opcode <= OPCODE_NOOP; -- When issuing an OPCODE, must be a pulse
    thrd2intrfc_address <= Z32;
    thrd2intrfc_value <= Z32;
    thrd2intrfc_function <= U_FUNCTION_USER_SELECT;
    next_state <= current_state;
    return_state_next <= return_state;

	arg_next <= arg;
	buffer_next <= bufer;
	bufLen_next <= bufLen;
	outputIndex_next <= outputIndex;
	index_next <= index;
	len_next <= len;
	pos_next <= pos;
	inputData_next <= inputData;
	outputData_next <= outputData;
	count_next <= count;

    -- The state machine
        case current_state is
          when FUNCTION_RESET =>
            --Set default values
            thrd2intrfc_opcode <= OPCODE_NOOP;
            thrd2intrfc_address <= Z32;
            thrd2intrfc_value <= Z32;
            thrd2intrfc_function <= U_FUNCTION_START;

			arg_next <= Z32;
			buffer_next <= Z32;
			bufLen_next <= Z32;
			outputIndex_next <= Z32;
			index_next <= Z32;
			len_next <= Z32;
			pos_next <= Z32;
			inputData_next <= Z32;
			outputData_next <= Z32;
			count_next <= Z32;

          when FUNCTION_START => 
            -- read the passed in argument
            thrd2intrfc_opcode <= OPCODE_POP;
            thrd2intrfc_address <= Z32;
            return_state_next <= READ_ARGS_1;
            next_state <= WAIT_STATE;
  
          -- int Code[MAX_SIZE]
          when READ_ARGS_1 =>
            arg_next <= toUser_value;
            -- Declare an array of MAX_SIZE on the stack
            thrd2intrfc_opcode <= OPCODE_DECLARE;
            thrd2intrfc_value <= MAX_SIZE;
            return_state_next <= READ_ARGS_2;
            next_state <= WAIT_STATE;

          -- struct HuffmanStructure * huffman = (struct HuffmanStructure *)arg;
          when READ_ARGS_2 =>
            -- Read value of inputData pointer
            thrd2intrfc_opcode <= OPCODE_LOAD;
            thrd2intrfc_address <= arg;
            return_state_next <= READ_ARGS_3;
            next_state <= WAIT_STATE;

          when READ_ARGS_3 => 
		    inputData_next <= toUser_value;
            -- Read value of outputData pointer
            thrd2intrfc_opcode <= OPCODE_LOAD;
            thrd2intrfc_address <= arg + 4;
            return_state_next <= READ_ARGS_4;
            next_state <= WAIT_STATE;

          when READ_ARGS_4 => 
		    outputData_next <= toUser_value;
            -- Read value of count
            thrd2intrfc_opcode <= OPCODE_LOAD;
            thrd2intrfc_address <= arg + 8;
            return_state_next <= READ_ARGS_5;
            next_state <= WAIT_STATE;

		  when READ_ARGS_5 =>
		    count_next <= toUser_value;
			next_state <= FORLOOP_1;

          -- for ( index = 0; index < huffman->count; index++ );
		  when FORLOOP_1 =>
		    -- index was initialized in the start state
			-- check to see if index is less than count
            if ( index < count ) then
			  next_state <= FORLOOP_2;
			else
			  next_state <= FLUSH_1;
			end if;

          -- Len = 0;
		  -- Pos = huffman->inputData[Index];
		  when FORLOOP_2 =>
		    -- len was initialized in the start state
			-- read the character to encode
            thrd2intrfc_opcode <= OPCODE_LOAD;
            thrd2intrfc_address <= inputData + (index(2 to 31) & "00");
            return_state_next <= FORLOOP_3;
            next_state <= WAIT_STATE;

		  when FORLOOP_3 =>
		    pos_next <= toUser_value;
			next_state <= WHILE_A_1;

          -- while ((pos < MAX_SIZE) && (huffman->code.Parent[Pos] >= 0 ))
		  when WHILE_A_1 =>
		    -- check to see if pos < MAX_SIZE
		    if ( pos < MAX_SIZE ) then
		      -- read the value of huffman->code.Parent[pos]
              thrd2intrfc_opcode <= OPCODE_LOAD;
              thrd2intrfc_address <= arg + x"0000100C" + (pos(2 to 31) & "00");
              return_state_next <= WHILE_A_2;
              next_state <= WAIT_STATE;
			else 
			  next_state <= WHILE_B_1;
			end if;

          -- code[len++] = huffman->code.bit[pos]
		  -- pos = huffman->code.parent[pos]
		  when WHILE_A_2 =>
		    -- check to see of huffman->code.Parent[pos] >= 0
			-- can check this by inspecting the bit 0
			case toUser_value(0) is
			  when '0' => 
			    -- this is a positive number or zero
                pos_next <= toUser_value;
		        -- read the value of huffman->code.bit[pos]
                thrd2intrfc_opcode <= OPCODE_LOAD;
                thrd2intrfc_address <= arg + x"0000400C" + (pos(2 to 31) & "00");
                return_state_next <= WHILE_A_3;
                next_state <= WAIT_STATE;
			  when others =>
			    -- this is a negative number
			    next_state <= WHILE_B_1;
			end case;

		  when WHILE_A_3 =>
		    -- set code[len] to the value of huffman->code.bit[pos]
		    thrd2intrfc_opcode <= OPCODE_WRITE;
			thrd2intrfc_value <= toUser_value;
			thrd2intrfc_address <= len;
			-- increment len
			len_next <= len + x"00000001";
			return_state_next <= WHILE_A_1;
			next_state <= WAIT_STATE;

		  -- end of while loop

          -- while( len > 0 )
		  when WHILE_B_1 =>
		    case len is
			  when x"00000000" =>
			    -- len is = 0
                next_state <= FORLOOP_4;
			  when others =>
			    -- len is > 0
				-- decrement len in preparation for next step
				len_next <= len - x"00000001";
				next_state <= WHILE_B_2;
			end case;

          -- Buffer = (Buffer << 1) | Code[--Len];
          when WHILE_B_2 =>
		    -- read the value of code[len]
		    thrd2intrfc_opcode <= OPCODE_READ;
			thrd2intrfc_value <= toUser_value;
			thrd2intrfc_address <= len;
			return_state_next <= WHILE_B_3;
			next_state <= WAIT_STATE;

          -- BufLen++;
		  when WHILE_B_3 =>
		    -- set the value of buffer
			--buffer_next <= (bufer(1 to 31) & '0') | toUser_value;
			buffer_next <= bufer(1 to 31) & toUser_value(31);
			-- increment buflen
			buflen_next <= bufLen + x"00000001";
			next_state <= WHILE_B_4;

		  -- if ( BufLen == 32 ) 
		  --   huffman->outputData[outputIndex] = Buffer
		  when WHILE_B_4 =>
		    -- check to see if BufLen == 32, do this by checking bit 26
            case bufLen(26) is
			  when '0' =>
			    -- bufLen is less than 32
				next_state <= WHILE_B_1;
			  when others =>
			    -- bufLen is 32
				-- store the value of outputData[outputIndex]
		        thrd2intrfc_opcode <= OPCODE_STORE;
			    thrd2intrfc_value <= bufer;
			    thrd2intrfc_address <= outputData + (outputIndex(2 to 31) & "00");
			    return_state_next <= WHILE_B_5;
			    next_state <= WAIT_STATE;
			end case;

		  -- outputIndex++;
		  -- Buffer = 0;
		  -- BufLen = 0;
		  when WHILE_B_5 =>
		    outputIndex_next <= outputIndex + x"00000001";
			buffer_next <= Z32;
			bufLen_next <= Z32;
			next_state <= WHILE_B_1;

		  -- end if statement
		  -- end while loop

		  when FORLOOP_4 =>
		    -- increment index
			index_next <= index + x"00000001";
			next_state <= FORLOOP_1;

		  -- end for loop

          -- if ( bufLen != 0 )
          --   Buffer = Buffer << (32 - BufLen)
          when FLUSH_1 =>
		    -- check to see if bufLen is equal to 0, only have to check last 6 bits
			-- if it is not 0, check the value to know how much to shift buffer
		    case bufLen(26 to 31) is
			  when "000000" =>
			    next_state <= EXIT_THREAD;
			  when "000001" =>
			    buffer_next <= bufer(31) & Z32(0 to 30);
			    next_state <= FLUSH_2;
			  when "000010" =>
			    buffer_next <= bufer(30 to 31) & Z32(0 to 29);
			    next_state <= FLUSH_2;
			  when "000011" =>
			    buffer_next <= bufer(29 to 31) & Z32(0 to 28);
			    next_state <= FLUSH_2;
			  when "000100" =>
			    buffer_next <= bufer(28 to 31) & Z32(0 to 27);
			    next_state <= FLUSH_2;
			  when "000101" =>
			    buffer_next <= bufer(27 to 31) & Z32(0 to 26);
			    next_state <= FLUSH_2;
			  when "000110" =>
			    buffer_next <= bufer(26 to 31) & Z32(0 to 25);
			    next_state <= FLUSH_2;
			  when "000111" =>
			    buffer_next <= bufer(25 to 31) & Z32(0 to 24);
			    next_state <= FLUSH_2;
			  when "001000" =>
			    buffer_next <= bufer(24 to 31) & Z32(0 to 23);
			    next_state <= FLUSH_2;
			  when "001001" =>
			    buffer_next <= bufer(23 to 31) & Z32(0 to 22);
			    next_state <= FLUSH_2;
			  when "001010" =>
			    buffer_next <= bufer(22 to 31) & Z32(0 to 21);
			    next_state <= FLUSH_2;
			  when "001011" =>
			    buffer_next <= bufer(21 to 31) & Z32(0 to 20);
			    next_state <= FLUSH_2;
			  when "001100" =>
			    buffer_next <= bufer(20 to 31) & Z32(0 to 19);
			    next_state <= FLUSH_2;
			  when "001101" =>
			    buffer_next <= bufer(19 to 31) & Z32(0 to 18);
			    next_state <= FLUSH_2;
			  when "001110" =>
			    buffer_next <= bufer(18 to 31) & Z32(0 to 17);
			    next_state <= FLUSH_2;
			  when "001111" =>
			    buffer_next <= bufer(17 to 31) & Z32(0 to 16);
			    next_state <= FLUSH_2;
			  when "010000" =>
			    buffer_next <= bufer(16 to 31) & Z32(0 to 15);
			    next_state <= FLUSH_2;
			  when "010001" =>
			    buffer_next <= bufer(15 to 31) & Z32(0 to 14);
			    next_state <= FLUSH_2;
			  when "010010" =>
			    buffer_next <= bufer(14 to 31) & Z32(0 to 13);
			    next_state <= FLUSH_2;
			  when "010011" =>
			    buffer_next <= bufer(13 to 31) & Z32(0 to 12);
			    next_state <= FLUSH_2;
			  when "010100" =>
			    buffer_next <= bufer(12 to 31) & Z32(0 to 11);
			    next_state <= FLUSH_2;
			  when "010101" =>
			    buffer_next <= bufer(11 to 31) & Z32(0 to 10);
			    next_state <= FLUSH_2;
			  when "010110" =>
			    buffer_next <= bufer(10 to 31) & Z32(0 to 9);
			    next_state <= FLUSH_2;
			  when "010111" =>
			    buffer_next <= bufer(9 to 31) & Z32(0 to 8);
			    next_state <= FLUSH_2;
			  when "011000" =>
			    buffer_next <= bufer(8 to 31) & Z32(0 to 7);
			    next_state <= FLUSH_2;
			  when "011001" =>
			    buffer_next <= bufer(7 to 31) & Z32(0 to 6);
			    next_state <= FLUSH_2;
			  when "011010" =>
			    buffer_next <= bufer(6 to 31) & Z32(0 to 5);
			    next_state <= FLUSH_2;
			  when "011011" =>
			    buffer_next <= bufer(5 to 31) & Z32(0 to 4);
			    next_state <= FLUSH_2;
			  when "011100" =>
			    buffer_next <= bufer(4 to 31) & Z32(0 to 3);
			    next_state <= FLUSH_2;
			  when "011101" =>
			    buffer_next <= bufer(3 to 31) & Z32(0 to 2);
			    next_state <= FLUSH_2;
			  when "011110" =>
			    buffer_next <= bufer(2 to 31) & Z32(0 to 1);
			    next_state <= FLUSH_2;
			  when "011111" =>
			    buffer_next <= bufer(1 to 31) & Z32(0);
			    next_state <= FLUSH_2;
			  when others =>
			    -- should never get to this state
			    next_state <= EXIT_THREAD;
		    end case;

		  -- huffman->outputData[outputIndex] = Buffer
		  when FLUSH_2 =>
		    thrd2intrfc_opcode <= OPCODE_STORE;
			thrd2intrfc_value <= bufer;
			thrd2intrfc_address <= outputData + (outputIndex(2 to 31) & "00");
			return_state_next <= EXIT_THREAD;
			next_state <= WAIT_STATE;

	      -- end if statement

          when EXIT_THREAD =>
		    thrd2intrfc_opcode <= OPCODE_PUSH;
			thrd2intrfc_value <= Z32;
			return_state_next <= EXIT_THREAD_1;
			next_state <= WAIT_STATE;

		  when EXIT_THREAD_1 =>
		    thrd2intrfc_opcode <= OPCODE_CALL;
			thrd2intrfc_value <= Z32;
			thrd2intrfc_function <= FUNCTION_HTHREAD_EXIT;
			next_state <= WAIT_STATE;

          when WAIT_STATE => 
            case toUser_goWait is
              when '1' => --Here because HWTUL chose to be here for one clock cycle
                next_state <= return_state;
              when OTHERS => --ie '0', Here because HWTI is telling us to wait
                next_state <= return_state;
            end case;

          when others =>
            next_state <= ERROR_STATE;

        end case;
      
  end process HWTUL_STATE_MACHINE;
end architecture IMP;
